// CSCB58 Winter 2017 Final Project
// Cave Catchers
// Names: Nathan Seebarran, Sadman Rafid, Kareem Hage-Ali, Raphael Ambegia 
// Description: Catch Yellows(+1)
//					 Catch Cyans(+5!)
//					 Avoid Reds(-10!!)
//					 gg

module GuitarBand
	(
		CLOCK_50,						//	On Board 50 MHz
		// Your inputs and outputs here
        KEY,
        SW,
		// The ports below are for the VGA output.  Do not change.
		VGA_CLK,   						//	VGA Clock
		VGA_HS,							//	VGA H_SYNC
		VGA_VS,							//	VGA V_SYNC
		VGA_BLANK_N,						//	VGA BLANK
		VGA_SYNC_N,						//	VGA SYNC
		VGA_R,   						//	VGA Red[9:0]
		VGA_G,	 						//	VGA Green[9:0]
		VGA_B,   						//	VGA Blue[9:0]
		HEX0, 
		HEX1
	);

	input			CLOCK_50;				//	50 MHz
	input   [9:0]   SW;
	input   [3:0]   KEY;

	// Declare your inputs and outputs here
	// Do not change the following outputs
	output			VGA_CLK;   				//	VGA Clock
	output			VGA_HS;					//	VGA H_SYNC
	output			VGA_VS;					//	VGA V_SYNC
	output			VGA_BLANK_N;				//	VGA BLANK
	output			VGA_SYNC_N;				//	VGA SYNC
	output	[9:0]	VGA_R;   				//	VGA Red[9:0]
	output	[9:0]	VGA_G;	 				//	VGA Green[9:0]
	output	[9:0]	VGA_B;   				//	VGA Blue[9:0]
	
	
	output [6:0] HEX0, HEX1;

	wire resetn;
	assign resetn = KEY[0];
	
	// Create the colour, x, y and writeEn wires that are inputs to the controller.
	wire [2:0] colour;
	wire [7:0] x;
	wire [6:0] y;
	wire writeEn;

	// Create an Instance of a VGA controller - there can be only one!
	// Define the number of colours as well as the initial ground
	// image file (.MIF) for the controller.
	vga_adapter VGA(
			.resetn(resetn),
			.clock(CLOCK_50),
			.colour(colour),
			.x(x),
			.y(y),
			.plot(1'b1),
			/* Signals for the DAC to drive the monitor. */
			.VGA_R(VGA_R),
			.VGA_G(VGA_G),
			.VGA_B(VGA_B),
			.VGA_HS(VGA_HS),
			.VGA_VS(VGA_VS),
			.VGA_BLANK(VGA_BLANK_N),
			.VGA_SYNC(VGA_SYNC_N),
			.VGA_CLK(VGA_CLK));
		defparam VGA.RESOLUTION = "160x120";
		defparam VGA.MONOCHROME = "FALSE";
		defparam VGA.BITS_PER_COLOUR_CHANNEL = 1;
		defparam VGA.BACKGROUND_IMAGE = "";
			
	// Put your code here. Your code should produce signals x,y,colour and writeEn/plot
	// for the VGA controller, in addition to any other functionality your design may require.
	wire [6:0] datain;
	wire load_x, load_y, load_r, load_c, ld_alu_out;
	wire go, loadEn;
	
	wire left, right;
	
	assign left = SW[2];
	assign right = SW[0];
	
	
	datapath d1(CLOCK_50, resetn, left, right, x, y, colour, data_result);

	
	wire [7:0] data_result;

	hex_decoder H0(
        .hex_digit(data_result[3:0]), 
        .segments(HEX0)
        );
        
    hex_decoder H1(
        .hex_digit(data_result[7:4]), 
        .segments(HEX1)
        );

    
endmodule

`define LANE_COUNT 2
`define LANE1_X 30
`define LANE2_X 90

`define HITBLOCK_Y 10

`define RED 3'b100
`define GREEN 3'b010
`define BLUE 3'b001
`define WHITE 3'b111
`define BLACK 3'b00

`define TICKS_PER_FRAME 500000


module datapath(
    input clk,
	 input resetn,
	 input left,
	 input right,
    output reg [7:0] x,
	 output reg [6:0] y,
	 output reg [2:0] colour,
	 output reg [7:0] data_result
    ); 
	 
	 
	//reg [4:0] ;
	reg pre_left;
	reg left_click;
	
	reg pre_right;
	reg right_click;
	
	reg [27:0] frame_counter;
	reg [3:0] lane_counter;
	reg [4:0] draw_counter;
	
    // output of the alu
   reg [7:0] x_alu;
	reg [6:0] y_alu;
	reg[4:0] count;
	reg[4:0] clear;
	reg[4:0] draw;
	
	// different falling blocks x and y registers

	reg [7:0] blockX1;
	reg [6:0] blockY1;
	reg [7:0] blockX2;
	reg [6:0] blockY2;
	
	initial begin 
		
		blockX1 <= `LANE1_X;
		blockY1 <= 0;
		blockX2 <= `LANE2_X;
		blockY2 <= 0;
		lane_counter <= 0;
		frame_counter <= 0;
		draw_counter <= 0;
		
		left_click <= 0;
		pre_left <= 1;
		right_click <= 0;
		pre_right <= 1;
	end
	
	
	
	always@(posedge clk) begin
		
		if(draw_counter == 2) begin
			draw_counter <= 0;
			// If we process every lane
			lane_counter <= lane_counter + 1;
			if(lane_counter == `LANE_COUNT) begin
				lane_counter <= 0;
				// Once every lane is proccesed, increment tick
				frame_counter <= frame_counter + 1;
				// If we reach the ticks per frame
				if(frame_counter == `TICKS_PER_FRAME) begin
					frame_counter <= 0;
				end
			end
		end

		
		// Update Lane 1
		if(lane_counter == 0) begin
			pre_left <= left;
			if(left == 1 && pre_left == 0) begin
				left_click <= 1;
			end
			if(draw_counter == 0 && left_click == 0) begin
				if (frame_counter == 0) begin
					x <= `LANE1_X;
					y <= `HITBLOCK_Y;
					colour <= `BLACK;
				end
			end
			if(draw_counter == 0 && left_click == 1) begin
				x <= `LANE1_X;
				y <= `HITBLOCK_Y;
				colour <= `WHITE;
				left_click <= 0;
			end
			if(draw_counter == 1) begin
				x <= blockX1;
				y <= blockY1;			
				colour <= `RED;
				if (frame_counter == 0) begin
					blockY1 <= blockY1 + 1;		
				end
			end
		end
		// Update Lane 2
		else if(lane_counter == 1) begin
			pre_right <= right;
			if(right == 1 && pre_right == 0) begin
				right_click <= 1;
			end
	
			if(draw_counter == 0 && right_click == 0) begin
				if (frame_counter == 0) begin
					x <= `LANE2_X;
					y <= `HITBLOCK_Y;
					colour <= `BLACK;
				end
			end
			else if(draw_counter == 0 && right_click == 1) begin
				x <= `LANE2_X;
				y <= `HITBLOCK_Y;
				colour <= `WHITE;
				right_click <= 0;
			end
			else if(draw_counter == 1) begin
				x <= blockX2;
				y <= blockY2;			
				colour <= `GREEN;
				if (frame_counter == 0) begin
					blockY2 <= blockY2 + 1;		
				end
			end
		end
		/*
		else if(lane_counter == 1) begin
			x <= blockX2;
			y <= blockY2;			
			colour <= `GREEN;
			if (frame_counter == 0) begin
				blockY2 <= blockY2 + 1;
			end	
		end
		*/
		// Go to next lane
		draw_counter <= draw_counter + 1;
	end

endmodule

// hex display
module hex_decoder(hex_digit, segments);
    input [3:0] hex_digit;
    output reg [6:0] segments;
   
    always @(*)
        case (hex_digit)
            4'h0: segments = 7'b100_0000;
            4'h1: segments = 7'b111_1001;
            4'h2: segments = 7'b010_0100;
            4'h3: segments = 7'b011_0000;
            4'h4: segments = 7'b001_1001;
            4'h5: segments = 7'b001_0010;
            4'h6: segments = 7'b000_0010;
            4'h7: segments = 7'b111_1000;
            4'h8: segments = 7'b000_0000;
            4'h9: segments = 7'b001_1000;
            4'hA: segments = 7'b000_1000;
            4'hB: segments = 7'b000_0011;
            4'hC: segments = 7'b100_0110;
            4'hD: segments = 7'b010_0001;
            4'hE: segments = 7'b000_0110;
            4'hF: segments = 7'b000_1110;   
            default: segments = 7'h7f;
        endcase
endmodule

